module top(input spiClk, input spiIn, output spiOut);

	assign spiOut = spiIn;

endmodule